----------------------------------------------------------------------------------
-- Company: EPFL
-- Engineer: Simon Thür
-- 
-- Create Date: 02.12.2022 22:27:12
-- Design Name: 
-- Module Name: pong_fsm_tb - Behavioral
-- Project Name: PONG
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------



library ieee;
library std;
-- Standard packages
use std.env.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- Packages
library work;
use work.dsd_prj_pkg.all;


entity pong_fsm_tb is
--  Port ( );
end pong_fsm_tb;

architecture Behavioral of pong_fsm_tb is

begin


end Behavioral;

thuer@DESKTOP-UUUA4G2.9120:1670770858
--=============================================================================
-- @file key_lock_timed.vhdl
-- @author Simon Thür
--=============================================================================
-- Standard library
library ieee;
-- Standard packages
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- =============================================================================

-- Keylock

-- @brief Keylock circuit for Lab3

-- =============================================================================